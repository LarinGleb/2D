break/192, 832/1;break/256, 832/1;break/512, 832/1;break/448, 832/1;break/448, 896/2;break/512, 896/2;break/576, 896/1;break/640, 896/1;
-1402,793
-30,8
393151
0:0:0;1:0:0;2:0:0;3:0:0;4:0:0;5:0:0;6:0:0;7:0:0;8:0:0;9:0:0;