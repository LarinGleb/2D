break/192, 832/1;break/256, 832/1;break/512, 832/1;break/448, 832/1;break/448, 896/2;break/512, 896/2;break/576, 896/1;break/640, 896/1;break/-1536, 896/1;break/-1472, 896/1;create/-1280, 768/1;create/-1280, 704/1;break/-1792, 896/1;break/-1728, 896/1;break/-1664, 896/1;break/-1600, 896/1;break/-1472, 960/2;break/-1472, 1024/3;break/-1536, 960/2;break/-1536, 1024/3;break/-1600, 960/2;break/-1600, 1024/3;break/-1664, 960/2;break/-1664, 1024/3;break/-1728, 960/2;break/-1728, 1024/3;break/-1792, 960/2;break/-1792, 1024/3;break/-1856, 960/1;create/-1664, 832/3;create/-1728, 896/3;create/-1792, 960/3;create/-1728, 704/3;create/-1600, 832/3;create/-1472, 896/3;create/-1984, 896/2;create/-1856, 832/2;create/-1856, 832/2;create/-2048, 704/2;create/-2048, 832/2;create/-1984, 896/2;
-2112,896
-46,8
393151
0:1:5;1:0:0;2:0:0;3:0:0;4:0:0;5:0:0;6:0:0;7:0:0;8:0:0;9:0:0;