break/-448, 768/1;break/-384, 768/1;break/-512, 768/1;break/-576, 768/1;create/-448, 576/1;create/-384, 640/1;create/-448, 704/1;create/-512, 640/1;break/-640, 896/2;break/-576, 832/2;break/-512, 832/2;break/-576, 896/3;break/-640, 832/1;break/-512, 896/3;break/-704, 832/1;create/-832, 576/3;create/-704, 640/3;create/-1472, 640/2;create/-1408, 704/2;create/-1408, 768/2;
-18966,5745
-302,8
429645
0:0:0;1:0:0;2:0:0;3:0:0;4:0:0;5:0:0;6:0:0;7:0:0;8:0:0;9:0:0;